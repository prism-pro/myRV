
//--xuezhen--

`include "defines.v"

module if_stage(
  input wire clk,
  input wire rst,
  input wire pc_op1,
  input wire pc_op2,
  input wire `REG_BUS rs1_data,
  input wire `REG_BUS imm_data,

  output wire `REG_BUS inst_addr,
  output wire         inst_ena
  
);

reg [`REG_BUS]pc;

// fetch an instruction
always@( posedge clk )
begin
  if( rst == 1'b1 )
  begin
    pc <= `ZERO_WORD ;
  end
  else
  begin
    pc <= pc + 4;
  end
end

assign inst_addr = pc;
assign inst_ena  = ( rst == 1'b1 ) ? 0 : 1;


endmodule
